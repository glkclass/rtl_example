`timescale 1ns/1ns
package dut_test_pkg;
    import uvm_pkg::*;
    `include "uvm_macros.svh"

    import typedef_pkg::*;
    import dut_tb_param_pkg::*;
    import dut_handler_pkg::*;
    import dut_env_pkg::*;
    import dut_agent_pkg::*;
    import dut_scb_pkg::*;
    import dut_sequence_pkg::*;
    `include "dut_test_base.svh"
    `include "dut_test.svh"
    `include "recorded_txn_test.svh"
endpackage




