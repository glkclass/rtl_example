`timescale 1ns/1ns
package dut_handler_pkg;
    import uvm_pkg::*;
    `include "uvm_macros.svh"

    import dut_tb_param_pkg::*;
    import typedef_pkg::*;
    `include "dut_report_server.svh"
    `include "dut_progress_bar.svh"
    `include "dut_handler.svh"
endpackage




