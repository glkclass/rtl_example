package typedef_pkg;
    typedef     int                     vector [];

    typedef     enum    {
                            IDLE = 0,
                            READ = 1,
                            WRITE = 2
                        }               t_recorder_db_mode;



endpackage

